----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:43:01 02/18/2015 
-- Design Name: 
-- Module Name:    RISCCONSTANTS_PKG - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package RISCCONSTANTS_PKG is
	constant DATAPATH		: integer := 16;		-- data width of RISC machine
end RISCCONSTANTS_PKG;

package body RISCCONSTANTS_PKG is

end RISCCONSTANTS_PKG;

