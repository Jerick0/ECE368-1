--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:21:21 03/24/2015
-- Design Name:   
-- Module Name:   C:/Users/Logan Doonan/Documents/Xilinx/ECE-368_Lab3/User_interface/tb_bank.vhd
-- Project Name:  User_interface
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: result_bank
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_bank IS
END tb_bank;
 
ARCHITECTURE behavior OF tb_bank IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT result_bank
    PORT(
         read_addr : IN  std_logic_vector(7 downto 0);
         data_in : IN  std_logic_vector(15 downto 0);
         data_out : OUT  std_logic_vector(15 downto 0);
         rst : IN  std_logic;
         w_en : IN  std_logic_vector(0 downto 0);
         clk : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal read_addr : std_logic_vector(7 downto 0) := (others => '0');
   signal data_in : std_logic_vector(15 downto 0) := (others => '0');
   signal rst : std_logic := '0';
   signal w_en : std_logic_vector(0 downto 0) := (others => '0');
   signal clk : std_logic := '0';

 	--Outputs
   signal data_out : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: result_bank PORT MAP (
          read_addr => read_addr,
          data_in => data_in,
          data_out => data_out,
          rst => rst,
          w_en => w_en,
          clk => clk
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		
      -- insert stimulus here 
		W_EN <= "1";
		wait for CLK_period;
		
		DATA_IN <= "0000000000000000";	--load instructions
		wait for CLK_period;
		DATA_IN <= "1111111111111111";	--load instructions
		wait for CLK_period;
		DATA_IN <= "0101010101010101";	--load instructions
		wait for CLK_period;
		DATA_IN <= "1010101010101010";	--load instructions
		wait for CLK_period*5;
		
		read_addr <= "00000001";	--load instructions
		wait for CLK_period;
		read_addr <= "00000010";	--load instructions
		wait for CLK_period;
		read_addr <= "00000011";	--load instructions
		wait for CLK_period;
		read_addr <= "00000100";	--load instructions

      wait;
   end process;

END;
